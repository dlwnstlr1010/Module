module big_mux_1bit (
    input [255:0] in, //1bit x 256 = 1024bit
    input [7:0] sel,
    output out);

    assign out = in[sel];
    
endmodule

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module big_1_mux_4bit (
    input [1023:0] in, //4bit x 256 = 1024bit
    input [7:0] sel,
    output [3:0] out);

    assign out = in[sel*4+:4]; // (sel*4) -> indexing, +:4 -> 4bit selecting
   
endmodule